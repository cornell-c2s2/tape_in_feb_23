VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO FFTSPIMinionRTL
  CLASS BLOCK ;
  FOREIGN FFTSPIMinionRTL ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 1760.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 0.000 700.030 4.000 ;
    END
  END clk
  PIN cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 146.920 2800.000 147.520 ;
    END
  END cs
  PIN cs_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 440.000 2800.000 440.600 ;
    END
  END cs_2
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END io_oeb[1]
  PIN miso
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1539.560 4.000 1540.160 ;
    END
  END miso
  PIN miso_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1099.600 4.000 1100.200 ;
    END
  END miso_2
  PIN mosi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 733.080 2800.000 733.680 ;
    END
  END mosi
  PIN mosi_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1026.160 2800.000 1026.760 ;
    END
  END mosi_2
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2099.530 0.000 2099.810 4.000 ;
    END
  END reset
  PIN sclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1319.240 2800.000 1319.840 ;
    END
  END sclk
  PIN sclk_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2796.000 1612.320 2800.000 1612.920 ;
    END
  END sclk_2
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2632.240 10.640 2633.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2785.840 10.640 2787.440 1749.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.040 10.640 2710.640 1749.200 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2794.040 1749.045 ;
      LAYER met1 ;
        RECT 5.520 10.640 2794.040 1749.200 ;
      LAYER met2 ;
        RECT 6.990 4.280 2788.430 1749.145 ;
        RECT 6.990 4.000 699.470 4.280 ;
        RECT 700.310 4.000 2099.250 4.280 ;
        RECT 2100.090 4.000 2788.430 4.280 ;
      LAYER met3 ;
        RECT 4.000 1613.320 2796.000 1749.125 ;
        RECT 4.000 1611.920 2795.600 1613.320 ;
        RECT 4.000 1540.560 2796.000 1611.920 ;
        RECT 4.400 1539.160 2796.000 1540.560 ;
        RECT 4.000 1320.240 2796.000 1539.160 ;
        RECT 4.000 1318.840 2795.600 1320.240 ;
        RECT 4.000 1100.600 2796.000 1318.840 ;
        RECT 4.400 1099.200 2796.000 1100.600 ;
        RECT 4.000 1027.160 2796.000 1099.200 ;
        RECT 4.000 1025.760 2795.600 1027.160 ;
        RECT 4.000 734.080 2796.000 1025.760 ;
        RECT 4.000 732.680 2795.600 734.080 ;
        RECT 4.000 660.640 2796.000 732.680 ;
        RECT 4.400 659.240 2796.000 660.640 ;
        RECT 4.000 441.000 2796.000 659.240 ;
        RECT 4.000 439.600 2795.600 441.000 ;
        RECT 4.000 220.680 2796.000 439.600 ;
        RECT 4.400 219.280 2796.000 220.680 ;
        RECT 4.000 147.920 2796.000 219.280 ;
        RECT 4.000 146.520 2795.600 147.920 ;
        RECT 4.000 10.715 2796.000 146.520 ;
      LAYER met4 ;
        RECT 822.775 558.455 865.440 1125.225 ;
        RECT 867.840 558.455 942.240 1125.225 ;
        RECT 944.640 558.455 1019.040 1125.225 ;
        RECT 1021.440 558.455 1095.840 1125.225 ;
        RECT 1098.240 558.455 1172.640 1125.225 ;
        RECT 1175.040 558.455 1249.440 1125.225 ;
        RECT 1251.840 558.455 1326.240 1125.225 ;
        RECT 1328.640 558.455 1403.040 1125.225 ;
        RECT 1405.440 558.455 1479.840 1125.225 ;
        RECT 1482.240 558.455 1556.640 1125.225 ;
        RECT 1559.040 558.455 1633.440 1125.225 ;
        RECT 1635.840 558.455 1710.240 1125.225 ;
        RECT 1712.640 558.455 1787.040 1125.225 ;
        RECT 1789.440 558.455 1863.840 1125.225 ;
        RECT 1866.240 558.455 1940.640 1125.225 ;
        RECT 1943.040 558.455 2017.440 1125.225 ;
        RECT 2019.840 558.455 2094.240 1125.225 ;
        RECT 2096.640 558.455 2171.040 1125.225 ;
        RECT 2173.440 558.455 2200.345 1125.225 ;
  END
END FFTSPIMinionRTL
END LIBRARY

